
module chip (input io_11_0_0, output io_11_0_1);

wire io_11_0_0;
assign io_11_0_1 = io_11_0_0;


endmodule

