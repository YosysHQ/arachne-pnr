
module chip (output io_11_0_0, input io_11_0_1);

wire io_11_0_0;
assign io_11_0_0 = io_11_0_1;


endmodule

