
module chip ();



endmodule

